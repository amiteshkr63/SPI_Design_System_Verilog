`define SPI_READY 1
`define SPI_BUSY 0

`define WORD_LENGTH 8

`define MODE_POL_PHS_00 'b00
`define MODE_POL_PHS_01 'b01
`define MODE_POL_PHS_10 'b10
`define MODE_POL_PHS_11 'b11

`define SPI_MODE MODE_POL_PHS_00

`define CLK_PER_HALF_BIT 2
`define PCKT_OK 0
`define PCKT_NOT_OK 1

`define DATA_VALID 1
`define DATA_INVALID 0

`define TOTAL_EDGE_COUNT 16

`define DISCONNECTED_FROM_SLAVE 1
`define CONNECTED_FROM_SLAVE 0